// `include "constants.v"

// module collision_detector(
//     input wire [9:0] player_x,    // Position of player x
//     input wire [9:0] player_y,    // Position of player y
//     input wire [9:0] car_x1, car_x2, car_x3, car_x4, // Car positions in x
//     output reg collision          // Indication of collision
// );



//     // Always block to detect collision
//     always @(*) begin
//         // Initialize collision to 0

//         // Verifying collision with car 1
        
//     end

// endmodule