// module frog(
//    input wire SW1,
//    input wire SW2,
//    input wire SW3,
//    input wire SW4,
// );
// endmodule